entity EntitiyName is
end entity;

architecture enitiyArch of EntityName is
begin
    process is
    begin
        -- code
    end process;
end architecture;
