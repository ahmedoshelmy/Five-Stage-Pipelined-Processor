LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
ENTITY MEMORY IS
    GENERIC (
        CACHE_WORD_WIDTH : INTEGER := 16;
        ADDRESS_BITS : INTEGER := 12
    );
    PORT (
        EN : IN STD_LOGIC;
        RST : IN STD_LOGIC;
        CLK : IN STD_LOGIC;
        MEMR : IN STD_LOGIC;
        MEMW : IN STD_LOGIC;
        ADDRESS_BUS : IN STD_LOGIC_VECTOR(ADDRESS_BITS - 1 DOWNTO 0);
        DATAIN : IN STD_LOGIC_VECTOR(CACHE_WORD_WIDTH DOWNTO 0);
        MEMOUT : OUT STD_LOGIC_VECTOR(CACHE_WORD_WIDTH - 1 DOWNTO 0));
END ENTITY MEMORY;

ARCHITECTURE ARCHMEMORY OF MEMORY IS
    TYPE MEMORYTYPE IS ARRAY((2 ** ADDRESS_BITS) - 1 DOWNTO 0) OF STD_LOGIC_VECTOR(CACHE_WORD_WIDTH - 1 DOWNTO 0);
    SIGNAL CACHE : MEMORYTYPE;
BEGIN
    PROCESS (CLK) BEGIN
        IF EN = '1' AND RISING_EDGE(CLK) THEN
            IF MEMR = '1' THEN
                MEMOUT <= CACHE(TO_INTEGER (unsigned(ADDRESS_BUS)));
            END IF;
            IF MEMW = '1' THEN
                CACHE(TO_INTEGER(unsigned(ADDRESS_BUS))) <= DATAIN;
            END IF;
        END IF;
        IF RST = '1' THEN
            CACHE <= (OTHERS => (OTHERS => '0'));
        END IF;
    END PROCESS;
END ARCHMEMORY;

-- TO_INTEGER here IS used TO convert STDLOGIC VECTOR TO INTEGER